--
-- Copyright: 2013, Technical University of Denmark, DTU Compute
-- Author: Martin Schoeberl (martin@jopdesign.com)
--         Rasmus Bo Soerensen (rasmus@rbscloud.dk)
-- License: Simplified BSD License
--

-- VHDL top level for Patmos in Chisel on Altera de2-115 board
--
-- Includes some 'magic' VHDL code to generate a reset after FPGA configuration.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity patmos_top is
  port(
    clk : in  std_logic;
    oLedsPins_led : out std_logic_vector(8 downto 0);
    iKeysPins_key : in std_logic_vector(3 downto 0);
    oUartPins_txd : out std_logic;
    iUartPins_rxd : in  std_logic;
    oSRAM_A : out std_logic_vector(19 downto 0);
    SRAM_DQ : inout std_logic_vector(15 downto 0);
    oSRAM_CE_N : out std_logic;
    oSRAM_OE_N : out std_logic;
    oSRAM_WE_N : out std_logic;
    oSRAM_LB_N : out std_logic;
    oSRAM_UB_N : out std_logic;
    oAudio_dacDat	: out std_logic;
    oAudio_dacLrc	: out std_logic;
    iAudio_adcDat	: in std_logic;
    oAudio_adcLrc	: out std_logic;
    ioAudio_sdat	: inout std_logic;
    oAudio_sclk	: out std_logic;
    oAudio_bclk	: out std_logic;
    oAudio_xclk	: out std_logic
    );
end entity patmos_top;

architecture rtl of patmos_top is
  component Patmos is
    port(
      clk             : in  std_logic;
      reset           : in  std_logic;

      io_comConf_M_Cmd        : out std_logic_vector(2 downto 0);
      io_comConf_M_Addr       : out std_logic_vector(31 downto 0);
      io_comConf_M_Data       : out std_logic_vector(31 downto 0);
      io_comConf_M_ByteEn     : out std_logic_vector(3 downto 0);
      io_comConf_M_RespAccept : out std_logic;
      io_comConf_S_Resp       : in std_logic_vector(1 downto 0);
      io_comConf_S_Data       : in std_logic_vector(31 downto 0);
      io_comConf_S_CmdAccept  : in std_logic;

      io_comSpm_M_Cmd         : out std_logic_vector(2 downto 0);
      io_comSpm_M_Addr        : out std_logic_vector(31 downto 0);
      io_comSpm_M_Data        : out std_logic_vector(31 downto 0);
      io_comSpm_M_ByteEn      : out std_logic_vector(3 downto 0);
      io_comSpm_S_Resp        : in std_logic_vector(1 downto 0);
      io_comSpm_S_Data        : in std_logic_vector(31 downto 0);

      io_cpuInfoPins_id   : in  std_logic_vector(31 downto 0);
      io_cpuInfoPins_cnt  : in  std_logic_vector(31 downto 0);
      io_ledsPins_led : out std_logic_vector(8 downto 0);
      io_keysPins_key : in  std_logic_vector(3 downto 0);
      io_uartPins_tx  : out std_logic;
      io_uartPins_rx  : in  std_logic;

      io_sramCtrlPins_ramOut_addr : out std_logic_vector(19 downto 0);
      io_sramCtrlPins_ramOut_doutEna : out std_logic;
      io_sramCtrlPins_ramIn_din : in std_logic_vector(15 downto 0);
      io_sramCtrlPins_ramOut_dout : out std_logic_vector(15 downto 0);
      io_sramCtrlPins_ramOut_nce : out std_logic;
      io_sramCtrlPins_ramOut_noe : out std_logic;
      io_sramCtrlPins_ramOut_nwe : out std_logic;
      io_sramCtrlPins_ramOut_nlb : out std_logic;
      io_sramCtrlPins_ramOut_nub : out std_logic;

      io_audioInterfacePins_dacDat	: out std_logic;
      io_audioInterfacePins_dacLrc	: out std_logic;
      io_audioInterfacePins_adcDat	: in std_logic;
      io_audioInterfacePins_adcLrc	: out std_logic;
      io_audioInterfacePins_sdIn		: in std_logic;
      io_audioInterfacePins_sdOut 	: out std_logic;
      io_audioInterfacePins_we 		: out std_logic;
      io_audioInterfacePins_sclkOut 	: out std_logic;
      io_audioInterfacePins_bclk		: out std_logic;
      io_audioInterfacePins_xclk		: out std_logic

      );
  end component;

  -- DE2-70: 50 MHz clock => 80 MHz
  -- BeMicro: 16 MHz clock => 25.6 MHz
  constant pll_infreq : real    := 50.0;
  constant pll_mult   : natural := 8;
  constant pll_div    : natural := 5;

  signal clk_int : std_logic;

  -- for generation of internal reset
  signal int_res            : std_logic;
  signal res_reg1, res_reg2 : std_logic;
  signal res_cnt            : unsigned(2 downto 0) := "000"; -- for the simulation

  -- sram signals for tristate inout
  signal sram_out_dout_ena : std_logic;
  signal sram_out_dout : std_logic_vector(15 downto 0);

  -- audio siganls for tristate inout
  signal saudio_sdIn		: std_logic;
  signal saudio_sdOut 	: std_logic;
  signal saudio_we 		: std_logic;
  signal saudio_sclkOut 	: std_logic;

  attribute altera_attribute : string;
  attribute altera_attribute of res_cnt : signal is "POWER_UP_LEVEL=LOW";

begin
  pll_inst : entity work.pll generic map(
    input_freq  => pll_infreq,
    multiply_by => pll_mult,
    divide_by   => pll_div
    )
    port map(
      inclk0 => clk,
      c0     => clk_int
      );
  -- we use a PLL
  -- clk_int <= clk;

  --
  --	internal reset generation
  --	should include the PLL lock signal
  --
  process(clk_int)
  begin
    if rising_edge(clk_int) then
      if (res_cnt /= "111") then
        res_cnt <= res_cnt + 1;
      end if;
      res_reg1 <= not res_cnt(0) or not res_cnt(1) or not res_cnt(2);
      res_reg2 <= res_reg1;
      int_res  <= res_reg2;
    end if;
  end process;


  -- tristate output to ssram
  process(sram_out_dout_ena, sram_out_dout)
  begin
    if sram_out_dout_ena='1' then
      SRAM_DQ <= sram_out_dout;
    else
      SRAM_DQ <= (others => 'Z');
    end if;
  end process;


  -- Audio I2C tristate buffer control
  --ioAudio_sdat <= saudio_sdOut when (saudio_we  = '0') else 'Z';
  --saudio_sdIn <= ioAudio_sdat when (saudio_we ='1') else '1';
  process(saudio_we, saudio_sdOut)
  begin
    if saudio_we = '1' then
      ioAudio_sdat <= saudio_sdOut;
      saudio_sdIn <= '1';
    else
      ioAudio_sdat <= 'Z';
      saudio_sdIn <= ioAudio_sdat;
    end if;
  end process;


  -- Not tristate
  oAudio_sclk <= saudio_sclkOut;

  comp : Patmos port map(clk_int, int_res,
                         open, open, open, open, open,
                         (others => '0'), (others => '0'), '0',
                         open, open, open, open,
                         (others => '0'), (others => '0'),
                         X"00000000", X"00000001",
                         oLedsPins_led,
                         iKeysPins_key,
                         oUartPins_txd, iUartPins_rxd,
                         oSRAM_A, sram_out_dout_ena, SRAM_DQ, sram_out_dout, oSRAM_CE_N, oSRAM_OE_N, oSRAM_WE_N, oSRAM_LB_N, oSRAM_UB_N,
                         oAudio_dacDat, oAudio_dacLrc, iAudio_adcDat, oAudio_adcLrc, saudio_sdIn, saudio_sdOut, saudio_we, saudio_sclkOut, oAudio_bclk, oAudio_xclk );

end architecture rtl;
