-- 
-- Copyright Technical University of Denmark. All rights reserved.
-- This file is part of the time-predictable VLIW Patmos.
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
-- 
--    1. Redistributions of source code must retain the above copyright notice,
--       this list of conditions and the following disclaimer.
-- 
--    2. Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDER ``AS IS'' AND ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES
-- OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN
-- NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF
-- THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation are
-- those of the authors and should not be interpreted as representing official
-- policies, either expressed or implied, of the copyright holder.
-- 


--------------------------------------------------------------------------------
-- Short descripton.
--
-- Author: Sahar Abbaspour
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity patmos_data_memory is
  generic (width : integer := 32; addr_width : integer := 10);
  port(
        clk       	             : in std_logic;
        wr_address               : in std_logic_vector(31 downto 0);
        data_in                  : in std_logic_vector(31 downto 0); -- store
        write_enable             : in std_logic;
        rd_address               : in std_logic_vector(31 downto 0);
        data_out                 : out std_logic_vector(31 downto 0) -- load
      );
end entity patmos_data_memory;

architecture arch of patmos_data_memory is
  -- TODO: define size and address range as a constant
  
  type data_memory is array (0 to 2**addr_width - 1) of std_logic_vector(width - 1 downto 0);
  signal data_mem : data_memory;

begin
  mem : process(clk)
  begin
  if (rising_edge(clk)) then
  	  data_out <= data_mem(to_integer(unsigned(rd_address(addr_width - 1 downto 0))));	
      if(write_enable = '1') then
        data_mem(to_integer(unsigned(wr_address(addr_width - 1 downto 0)))) <= data_in;
      end if;
    end if;
  end process mem;
end arch;
